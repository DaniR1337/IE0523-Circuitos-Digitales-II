module RX(  input   CKP, CPH, SCK, SS, MOSI,
            output  MISO);

endmodule
