module atm(CLK, RESET, TARJETA_RECIBIDA, PIN, DIGITO, DIGITO_STB, TIPO_TRANS, MONTO, MONTO_STB, BALANCE_ACTUALIZADO, ENTREGAR_DINERO, FONDOS_INSUFICIENTES, PIN_INCORRECTO, ADVERTENCIA, BLOQUEO);

// Inputs
input  CLK, RESET, TARJETA_RECIBIDA, TIPO_TRANS, DIGITO_STB, MONTO_STB;
input [3:0] DIGITO;
input [15:0] PIN;
input [31:0] MONTO;

// Outputs
output ENTREGAR_DINERO, PIN_INCORRECTO, ADVERTENCIA, BLOQUEO, FONDOS_INSUFICIENTES, BALANCE_ACTUALIZADO;

// Registros interno
reg BALANCE, ESTADO, PROX_ESTADO;

// Descripción de Flip FLops
always @(posedge CLK) begin
    if (RESET) begin
        ESTADO <= 0;
    end else begin
        ESTADO <= PROX_ESTADO;
    end
end


endmodule
